library verilog;
use verilog.vl_types.all;
entity SpecialTestBench is
end SpecialTestBench;
