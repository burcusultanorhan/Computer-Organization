module SelectALUSource();

endmodule