library verilog;
use verilog.vl_types.all;
entity MIPS is
    port(
        clock           : in     vl_logic
    );
end MIPS;
