module _32bit_and(A,B,F);
	input [31:0] A,B;
	output [31:0] F;

	and g31(F[31],A[31],B[31]);
	and g30(F[30],A[30],B[30]);
	and g29(F[29],A[29],B[29]);	
	and g28(F[28],A[28],B[28]);
	and g27(F[27],A[27],B[27]);
	and g26(F[26],A[26],B[26]);
	and g25(F[25],A[25],B[25]);	
	and g24(F[24],A[24],B[24]);
	and g23(F[23],A[23],B[23]);
	and g22(F[22],A[22],B[22]);
	and g21(F[21],A[21],B[21]);	
	and g20(F[20],A[20],B[20]);
	and g19(F[19],A[19],B[19]);
	and g18(F[18],A[18],B[18]);
	and g17(F[17],A[17],B[17]);	
	and g16(F[16],A[16],B[16]);
	and g15(F[15],A[15],B[15]);
	and g14(F[14],A[14],B[14]);
	and g13(F[13],A[13],B[13]);	
	and g12(F[12],A[12],B[12]);
	and g11(F[11],A[11],B[11]);
	and g10(F[10],A[10],B[10]);
	and g9(F[9],A[9],B[9]);	
	and g8(F[8],A[8],B[8]);
	and g7(F[7],A[7],B[7]);
	and g6(F[6],A[6],B[6]);
	and g5(F[5],A[5],B[5]);	
	and g4(F[4],A[4],B[4]);
	and g3(F[3],A[3],B[3]);
	and g2(F[2],A[2],B[2]);
	and g1(F[1],A[1],B[1]);	
	and g0(F[0],A[0],B[0]);
	
endmodule