library verilog;
use verilog.vl_types.all;
entity MIPS_testbench is
end MIPS_testbench;
